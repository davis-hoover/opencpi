../adc_samp_drop_generator/data_src.vhd