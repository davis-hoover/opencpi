../cdc_bits_tester.hdl/mmcm_100_to_100_50_and_25_top.vhd