../cdc_bits_tester.hdl/cdc_clk_gen.vhd