../../../../platform/hdl/primitives/zynq_ultra/zynq_ultra_pkg.vhd