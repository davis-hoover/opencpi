../data_sink_qdac_ad9361_sub.hdl/clock_selector_with_async_select.vhd