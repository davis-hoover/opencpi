../data_sink_qdac_ad9361_sub.hdl/clock_divider.vhd