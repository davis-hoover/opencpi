../time_corrector/file_writer.vhd