../adc_samp_drop_detector/data_src.vhd