../cdc_bits_tester.hdl/gen_clk.vhd