../event_in_x2_to_txen_tester.hdl/event_in_to_txen.vhd