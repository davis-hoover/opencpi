../adc_samp_drop_generator/file_writer.vhd