../../../../platform/hdl/primitives/zynq/zynq_pkg.vhd