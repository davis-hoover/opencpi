../rfdc_adc_config_0.hdl/rfdc_adc_config_0.vhd