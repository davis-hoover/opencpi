../../../../assets/hdl/devices/ad9361_dac_sub.hdl/event_in_x2_to_txen.vhd