../adc_samp_drop_detector/file_writer.vhd